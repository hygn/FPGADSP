module lut ( input en, input[6:0] lookup, output[7:0] out);
always @(en)begin
    case (lookup)
        7'd0: out <= 8'd127;
        7'd1: out <= 8'd133;
        7'd2: out <= 8'd140;
        7'd3: out <= 8'd146;
        7'd4: out <= 8'd152;
        7'd5: out <= 8'd158;
        7'd6: out <= 8'd164;
        7'd7: out <= 8'd170;
        7'd8: out <= 8'd176;
        7'd9: out <= 8'd182;
        7'd10: out <= 8'd187;
        7'd11: out <= 8'd193;
        7'd12: out <= 8'd198;
        7'd13: out <= 8'd203;
        7'd14: out <= 8'd208;
        7'd15: out <= 8'd213;
        7'd16: out <= 8'd217;
        7'd17: out <= 8'd222;
        7'd18: out <= 8'd226;
        7'd19: out <= 8'd230;
        7'd20: out <= 8'd233;
        7'd21: out <= 8'd236;
        7'd22: out <= 8'd240;
        7'd23: out <= 8'd242;
        7'd24: out <= 8'd245;
        7'd25: out <= 8'd247;
        7'd26: out <= 8'd249;
        7'd27: out <= 8'd251;
        7'd28: out <= 8'd252;
        7'd29: out <= 8'd253;
        7'd30: out <= 8'd254;
        7'd31: out <= 8'd254;
        7'd32: out <= 8'd254;
        7'd33: out <= 8'd254;
        7'd34: out <= 8'd253;
        7'd35: out <= 8'd252;
        7'd36: out <= 8'd251;
        7'd37: out <= 8'd250;
        7'd38: out <= 8'd248;
        7'd39: out <= 8'd246;
        7'd40: out <= 8'd244;
        7'd41: out <= 8'd241;
        7'd42: out <= 8'd238;
        7'd43: out <= 8'd235;
        7'd44: out <= 8'd231;
        7'd45: out <= 8'd228;
        7'd46: out <= 8'd224;
        7'd47: out <= 8'd220;
        7'd48: out <= 8'd215;
        7'd49: out <= 8'd210;
        7'd50: out <= 8'd206;
        7'd51: out <= 8'd201;
        7'd52: out <= 8'd195;
        7'd53: out <= 8'd190;
        7'd54: out <= 8'd185;
        7'd55: out <= 8'd179;
        7'd56: out <= 8'd173;
        7'd57: out <= 8'd167;
        7'd58: out <= 8'd161;
        7'd59: out <= 8'd155;
        7'd60: out <= 8'd149;
        7'd61: out <= 8'd143;
        7'd62: out <= 8'd136;
        7'd63: out <= 8'd130;
        7'd64: out <= 8'd124;
        7'd65: out <= 8'd118;
        7'd66: out <= 8'd111;
        7'd67: out <= 8'd105;
        7'd68: out <= 8'd99;
        7'd69: out <= 8'd93;
        7'd70: out <= 8'd87;
        7'd71: out <= 8'd81;
        7'd72: out <= 8'd75;
        7'd73: out <= 8'd69;
        7'd74: out <= 8'd64;
        7'd75: out <= 8'd59;
        7'd76: out <= 8'd53;
        7'd77: out <= 8'd48;
        7'd78: out <= 8'd44;
        7'd79: out <= 8'd39;
        7'd80: out <= 8'd34;
        7'd81: out <= 8'd30;
        7'd82: out <= 8'd26;
        7'd83: out <= 8'd23;
        7'd84: out <= 8'd19;
        7'd85: out <= 8'd16;
        7'd86: out <= 8'd13;
        7'd87: out <= 8'd10;
        7'd88: out <= 8'd8;
        7'd89: out <= 8'd6;
        7'd90: out <= 8'd4;
        7'd91: out <= 8'd3;
        7'd92: out <= 8'd2;
        7'd93: out <= 8'd1;
        7'd94: out <= 8'd0;
        7'd95: out <= 8'd0;
        7'd96: out <= 8'd0;
        7'd97: out <= 8'd0;
        7'd98: out <= 8'd1;
        7'd99: out <= 8'd2;
        7'd100: out <= 8'd3;
        7'd101: out <= 8'd5;
        7'd102: out <= 8'd7;
        7'd103: out <= 8'd9;
        7'd104: out <= 8'd12;
        7'd105: out <= 8'd14;
        7'd106: out <= 8'd18;
        7'd107: out <= 8'd21;
        7'd108: out <= 8'd24;
        7'd109: out <= 8'd28;
        7'd110: out <= 8'd32;
        7'd111: out <= 8'd37;
        7'd112: out <= 8'd41;
        7'd113: out <= 8'd46;
        7'd114: out <= 8'd51;
        7'd115: out <= 8'd56;
        7'd116: out <= 8'd61;
        7'd117: out <= 8'd67;
        7'd118: out <= 8'd72;
        7'd119: out <= 8'd78;
        7'd120: out <= 8'd84;
        7'd121: out <= 8'd90;
        7'd122: out <= 8'd96;
        7'd123: out <= 8'd102;
        7'd124: out <= 8'd108;
        7'd125: out <= 8'd114;
        7'd126: out <= 8'd121;
        7'd127: out <= 8'd127;
    endcase
end
endmodule
