module lut ( input clk, input[9:0] lookup, output[7:0] sine);
always @(posedge clk)begin
    case (lookup)
        10'd0: sine <= 8'd127;
        10'd1: sine <= 8'd128;
        10'd2: sine <= 8'd129;
        10'd3: sine <= 8'd129;
        10'd4: sine <= 8'd130;
        10'd5: sine <= 8'd131;
        10'd6: sine <= 8'd132;
        10'd7: sine <= 8'd132;
        10'd8: sine <= 8'd133;
        10'd9: sine <= 8'd134;
        10'd10: sine <= 8'd135;
        10'd11: sine <= 8'd136;
        10'd12: sine <= 8'd136;
        10'd13: sine <= 8'd137;
        10'd14: sine <= 8'd138;
        10'd15: sine <= 8'd139;
        10'd16: sine <= 8'd139;
        10'd17: sine <= 8'd140;
        10'd18: sine <= 8'd141;
        10'd19: sine <= 8'd142;
        10'd20: sine <= 8'd143;
        10'd21: sine <= 8'd143;
        10'd22: sine <= 8'd144;
        10'd23: sine <= 8'd145;
        10'd24: sine <= 8'd146;
        10'd25: sine <= 8'd146;
        10'd26: sine <= 8'd147;
        10'd27: sine <= 8'd148;
        10'd28: sine <= 8'd149;
        10'd29: sine <= 8'd150;
        10'd30: sine <= 8'd150;
        10'd31: sine <= 8'd151;
        10'd32: sine <= 8'd152;
        10'd33: sine <= 8'd153;
        10'd34: sine <= 8'd153;
        10'd35: sine <= 8'd154;
        10'd36: sine <= 8'd155;
        10'd37: sine <= 8'd156;
        10'd38: sine <= 8'd156;
        10'd39: sine <= 8'd157;
        10'd40: sine <= 8'd158;
        10'd41: sine <= 8'd159;
        10'd42: sine <= 8'd159;
        10'd43: sine <= 8'd160;
        10'd44: sine <= 8'd161;
        10'd45: sine <= 8'd162;
        10'd46: sine <= 8'd162;
        10'd47: sine <= 8'd163;
        10'd48: sine <= 8'd164;
        10'd49: sine <= 8'd165;
        10'd50: sine <= 8'd165;
        10'd51: sine <= 8'd166;
        10'd52: sine <= 8'd167;
        10'd53: sine <= 8'd168;
        10'd54: sine <= 8'd168;
        10'd55: sine <= 8'd169;
        10'd56: sine <= 8'd170;
        10'd57: sine <= 8'd171;
        10'd58: sine <= 8'd171;
        10'd59: sine <= 8'd172;
        10'd60: sine <= 8'd173;
        10'd61: sine <= 8'd173;
        10'd62: sine <= 8'd174;
        10'd63: sine <= 8'd175;
        10'd64: sine <= 8'd176;
        10'd65: sine <= 8'd176;
        10'd66: sine <= 8'd177;
        10'd67: sine <= 8'd178;
        10'd68: sine <= 8'd179;
        10'd69: sine <= 8'd179;
        10'd70: sine <= 8'd180;
        10'd71: sine <= 8'd181;
        10'd72: sine <= 8'd181;
        10'd73: sine <= 8'd182;
        10'd74: sine <= 8'd183;
        10'd75: sine <= 8'd183;
        10'd76: sine <= 8'd184;
        10'd77: sine <= 8'd185;
        10'd78: sine <= 8'd186;
        10'd79: sine <= 8'd186;
        10'd80: sine <= 8'd187;
        10'd81: sine <= 8'd188;
        10'd82: sine <= 8'd188;
        10'd83: sine <= 8'd189;
        10'd84: sine <= 8'd190;
        10'd85: sine <= 8'd190;
        10'd86: sine <= 8'd191;
        10'd87: sine <= 8'd192;
        10'd88: sine <= 8'd192;
        10'd89: sine <= 8'd193;
        10'd90: sine <= 8'd194;
        10'd91: sine <= 8'd194;
        10'd92: sine <= 8'd195;
        10'd93: sine <= 8'd196;
        10'd94: sine <= 8'd196;
        10'd95: sine <= 8'd197;
        10'd96: sine <= 8'd198;
        10'd97: sine <= 8'd198;
        10'd98: sine <= 8'd199;
        10'd99: sine <= 8'd200;
        10'd100: sine <= 8'd200;
        10'd101: sine <= 8'd201;
        10'd102: sine <= 8'd201;
        10'd103: sine <= 8'd202;
        10'd104: sine <= 8'd203;
        10'd105: sine <= 8'd203;
        10'd106: sine <= 8'd204;
        10'd107: sine <= 8'd205;
        10'd108: sine <= 8'd205;
        10'd109: sine <= 8'd206;
        10'd110: sine <= 8'd206;
        10'd111: sine <= 8'd207;
        10'd112: sine <= 8'd208;
        10'd113: sine <= 8'd208;
        10'd114: sine <= 8'd209;
        10'd115: sine <= 8'd209;
        10'd116: sine <= 8'd210;
        10'd117: sine <= 8'd211;
        10'd118: sine <= 8'd211;
        10'd119: sine <= 8'd212;
        10'd120: sine <= 8'd212;
        10'd121: sine <= 8'd213;
        10'd122: sine <= 8'd214;
        10'd123: sine <= 8'd214;
        10'd124: sine <= 8'd215;
        10'd125: sine <= 8'd215;
        10'd126: sine <= 8'd216;
        10'd127: sine <= 8'd216;
        10'd128: sine <= 8'd217;
        10'd129: sine <= 8'd217;
        10'd130: sine <= 8'd218;
        10'd131: sine <= 8'd219;
        10'd132: sine <= 8'd219;
        10'd133: sine <= 8'd220;
        10'd134: sine <= 8'd220;
        10'd135: sine <= 8'd221;
        10'd136: sine <= 8'd221;
        10'd137: sine <= 8'd222;
        10'd138: sine <= 8'd222;
        10'd139: sine <= 8'd223;
        10'd140: sine <= 8'd223;
        10'd141: sine <= 8'd224;
        10'd142: sine <= 8'd224;
        10'd143: sine <= 8'd225;
        10'd144: sine <= 8'd225;
        10'd145: sine <= 8'd226;
        10'd146: sine <= 8'd226;
        10'd147: sine <= 8'd227;
        10'd148: sine <= 8'd227;
        10'd149: sine <= 8'd228;
        10'd150: sine <= 8'd228;
        10'd151: sine <= 8'd229;
        10'd152: sine <= 8'd229;
        10'd153: sine <= 8'd230;
        10'd154: sine <= 8'd230;
        10'd155: sine <= 8'd230;
        10'd156: sine <= 8'd231;
        10'd157: sine <= 8'd231;
        10'd158: sine <= 8'd232;
        10'd159: sine <= 8'd232;
        10'd160: sine <= 8'd233;
        10'd161: sine <= 8'd233;
        10'd162: sine <= 8'd234;
        10'd163: sine <= 8'd234;
        10'd164: sine <= 8'd234;
        10'd165: sine <= 8'd235;
        10'd166: sine <= 8'd235;
        10'd167: sine <= 8'd236;
        10'd168: sine <= 8'd236;
        10'd169: sine <= 8'd236;
        10'd170: sine <= 8'd237;
        10'd171: sine <= 8'd237;
        10'd172: sine <= 8'd238;
        10'd173: sine <= 8'd238;
        10'd174: sine <= 8'd238;
        10'd175: sine <= 8'd239;
        10'd176: sine <= 8'd239;
        10'd177: sine <= 8'd239;
        10'd178: sine <= 8'd240;
        10'd179: sine <= 8'd240;
        10'd180: sine <= 8'd241;
        10'd181: sine <= 8'd241;
        10'd182: sine <= 8'd241;
        10'd183: sine <= 8'd242;
        10'd184: sine <= 8'd242;
        10'd185: sine <= 8'd242;
        10'd186: sine <= 8'd243;
        10'd187: sine <= 8'd243;
        10'd188: sine <= 8'd243;
        10'd189: sine <= 8'd243;
        10'd190: sine <= 8'd244;
        10'd191: sine <= 8'd244;
        10'd192: sine <= 8'd244;
        10'd193: sine <= 8'd245;
        10'd194: sine <= 8'd245;
        10'd195: sine <= 8'd245;
        10'd196: sine <= 8'd246;
        10'd197: sine <= 8'd246;
        10'd198: sine <= 8'd246;
        10'd199: sine <= 8'd246;
        10'd200: sine <= 8'd247;
        10'd201: sine <= 8'd247;
        10'd202: sine <= 8'd247;
        10'd203: sine <= 8'd247;
        10'd204: sine <= 8'd248;
        10'd205: sine <= 8'd248;
        10'd206: sine <= 8'd248;
        10'd207: sine <= 8'd248;
        10'd208: sine <= 8'd249;
        10'd209: sine <= 8'd249;
        10'd210: sine <= 8'd249;
        10'd211: sine <= 8'd249;
        10'd212: sine <= 8'd249;
        10'd213: sine <= 8'd250;
        10'd214: sine <= 8'd250;
        10'd215: sine <= 8'd250;
        10'd216: sine <= 8'd250;
        10'd217: sine <= 8'd250;
        10'd218: sine <= 8'd251;
        10'd219: sine <= 8'd251;
        10'd220: sine <= 8'd251;
        10'd221: sine <= 8'd251;
        10'd222: sine <= 8'd251;
        10'd223: sine <= 8'd251;
        10'd224: sine <= 8'd252;
        10'd225: sine <= 8'd252;
        10'd226: sine <= 8'd252;
        10'd227: sine <= 8'd252;
        10'd228: sine <= 8'd252;
        10'd229: sine <= 8'd252;
        10'd230: sine <= 8'd252;
        10'd231: sine <= 8'd253;
        10'd232: sine <= 8'd253;
        10'd233: sine <= 8'd253;
        10'd234: sine <= 8'd253;
        10'd235: sine <= 8'd253;
        10'd236: sine <= 8'd253;
        10'd237: sine <= 8'd253;
        10'd238: sine <= 8'd253;
        10'd239: sine <= 8'd253;
        10'd240: sine <= 8'd253;
        10'd241: sine <= 8'd253;
        10'd242: sine <= 8'd254;
        10'd243: sine <= 8'd254;
        10'd244: sine <= 8'd254;
        10'd245: sine <= 8'd254;
        10'd246: sine <= 8'd254;
        10'd247: sine <= 8'd254;
        10'd248: sine <= 8'd254;
        10'd249: sine <= 8'd254;
        10'd250: sine <= 8'd254;
        10'd251: sine <= 8'd254;
        10'd252: sine <= 8'd254;
        10'd253: sine <= 8'd254;
        10'd254: sine <= 8'd254;
        10'd255: sine <= 8'd254;
        10'd256: sine <= 8'd254;
        10'd257: sine <= 8'd254;
        10'd258: sine <= 8'd254;
        10'd259: sine <= 8'd254;
        10'd260: sine <= 8'd254;
        10'd261: sine <= 8'd254;
        10'd262: sine <= 8'd254;
        10'd263: sine <= 8'd254;
        10'd264: sine <= 8'd254;
        10'd265: sine <= 8'd254;
        10'd266: sine <= 8'd254;
        10'd267: sine <= 8'd254;
        10'd268: sine <= 8'd254;
        10'd269: sine <= 8'd254;
        10'd270: sine <= 8'd254;
        10'd271: sine <= 8'd253;
        10'd272: sine <= 8'd253;
        10'd273: sine <= 8'd253;
        10'd274: sine <= 8'd253;
        10'd275: sine <= 8'd253;
        10'd276: sine <= 8'd253;
        10'd277: sine <= 8'd253;
        10'd278: sine <= 8'd253;
        10'd279: sine <= 8'd253;
        10'd280: sine <= 8'd253;
        10'd281: sine <= 8'd252;
        10'd282: sine <= 8'd252;
        10'd283: sine <= 8'd252;
        10'd284: sine <= 8'd252;
        10'd285: sine <= 8'd252;
        10'd286: sine <= 8'd252;
        10'd287: sine <= 8'd252;
        10'd288: sine <= 8'd252;
        10'd289: sine <= 8'd251;
        10'd290: sine <= 8'd251;
        10'd291: sine <= 8'd251;
        10'd292: sine <= 8'd251;
        10'd293: sine <= 8'd251;
        10'd294: sine <= 8'd251;
        10'd295: sine <= 8'd250;
        10'd296: sine <= 8'd250;
        10'd297: sine <= 8'd250;
        10'd298: sine <= 8'd250;
        10'd299: sine <= 8'd250;
        10'd300: sine <= 8'd249;
        10'd301: sine <= 8'd249;
        10'd302: sine <= 8'd249;
        10'd303: sine <= 8'd249;
        10'd304: sine <= 8'd248;
        10'd305: sine <= 8'd248;
        10'd306: sine <= 8'd248;
        10'd307: sine <= 8'd248;
        10'd308: sine <= 8'd248;
        10'd309: sine <= 8'd247;
        10'd310: sine <= 8'd247;
        10'd311: sine <= 8'd247;
        10'd312: sine <= 8'd246;
        10'd313: sine <= 8'd246;
        10'd314: sine <= 8'd246;
        10'd315: sine <= 8'd246;
        10'd316: sine <= 8'd245;
        10'd317: sine <= 8'd245;
        10'd318: sine <= 8'd245;
        10'd319: sine <= 8'd245;
        10'd320: sine <= 8'd244;
        10'd321: sine <= 8'd244;
        10'd322: sine <= 8'd244;
        10'd323: sine <= 8'd243;
        10'd324: sine <= 8'd243;
        10'd325: sine <= 8'd243;
        10'd326: sine <= 8'd242;
        10'd327: sine <= 8'd242;
        10'd328: sine <= 8'd242;
        10'd329: sine <= 8'd241;
        10'd330: sine <= 8'd241;
        10'd331: sine <= 8'd241;
        10'd332: sine <= 8'd240;
        10'd333: sine <= 8'd240;
        10'd334: sine <= 8'd240;
        10'd335: sine <= 8'd239;
        10'd336: sine <= 8'd239;
        10'd337: sine <= 8'd239;
        10'd338: sine <= 8'd238;
        10'd339: sine <= 8'd238;
        10'd340: sine <= 8'd237;
        10'd341: sine <= 8'd237;
        10'd342: sine <= 8'd237;
        10'd343: sine <= 8'd236;
        10'd344: sine <= 8'd236;
        10'd345: sine <= 8'd235;
        10'd346: sine <= 8'd235;
        10'd347: sine <= 8'd235;
        10'd348: sine <= 8'd234;
        10'd349: sine <= 8'd234;
        10'd350: sine <= 8'd233;
        10'd351: sine <= 8'd233;
        10'd352: sine <= 8'd232;
        10'd353: sine <= 8'd232;
        10'd354: sine <= 8'd232;
        10'd355: sine <= 8'd231;
        10'd356: sine <= 8'd231;
        10'd357: sine <= 8'd230;
        10'd358: sine <= 8'd230;
        10'd359: sine <= 8'd229;
        10'd360: sine <= 8'd229;
        10'd361: sine <= 8'd228;
        10'd362: sine <= 8'd228;
        10'd363: sine <= 8'd227;
        10'd364: sine <= 8'd227;
        10'd365: sine <= 8'd226;
        10'd366: sine <= 8'd226;
        10'd367: sine <= 8'd225;
        10'd368: sine <= 8'd225;
        10'd369: sine <= 8'd224;
        10'd370: sine <= 8'd224;
        10'd371: sine <= 8'd223;
        10'd372: sine <= 8'd223;
        10'd373: sine <= 8'd222;
        10'd374: sine <= 8'd222;
        10'd375: sine <= 8'd221;
        10'd376: sine <= 8'd221;
        10'd377: sine <= 8'd220;
        10'd378: sine <= 8'd220;
        10'd379: sine <= 8'd219;
        10'd380: sine <= 8'd219;
        10'd381: sine <= 8'd218;
        10'd382: sine <= 8'd218;
        10'd383: sine <= 8'd217;
        10'd384: sine <= 8'd217;
        10'd385: sine <= 8'd216;
        10'd386: sine <= 8'd215;
        10'd387: sine <= 8'd215;
        10'd388: sine <= 8'd214;
        10'd389: sine <= 8'd214;
        10'd390: sine <= 8'd213;
        10'd391: sine <= 8'd213;
        10'd392: sine <= 8'd212;
        10'd393: sine <= 8'd211;
        10'd394: sine <= 8'd211;
        10'd395: sine <= 8'd210;
        10'd396: sine <= 8'd210;
        10'd397: sine <= 8'd209;
        10'd398: sine <= 8'd209;
        10'd399: sine <= 8'd208;
        10'd400: sine <= 8'd207;
        10'd401: sine <= 8'd207;
        10'd402: sine <= 8'd206;
        10'd403: sine <= 8'd206;
        10'd404: sine <= 8'd205;
        10'd405: sine <= 8'd204;
        10'd406: sine <= 8'd204;
        10'd407: sine <= 8'd203;
        10'd408: sine <= 8'd202;
        10'd409: sine <= 8'd202;
        10'd410: sine <= 8'd201;
        10'd411: sine <= 8'd201;
        10'd412: sine <= 8'd200;
        10'd413: sine <= 8'd199;
        10'd414: sine <= 8'd199;
        10'd415: sine <= 8'd198;
        10'd416: sine <= 8'd197;
        10'd417: sine <= 8'd197;
        10'd418: sine <= 8'd196;
        10'd419: sine <= 8'd195;
        10'd420: sine <= 8'd195;
        10'd421: sine <= 8'd194;
        10'd422: sine <= 8'd193;
        10'd423: sine <= 8'd193;
        10'd424: sine <= 8'd192;
        10'd425: sine <= 8'd191;
        10'd426: sine <= 8'd191;
        10'd427: sine <= 8'd190;
        10'd428: sine <= 8'd189;
        10'd429: sine <= 8'd189;
        10'd430: sine <= 8'd188;
        10'd431: sine <= 8'd187;
        10'd432: sine <= 8'd187;
        10'd433: sine <= 8'd186;
        10'd434: sine <= 8'd185;
        10'd435: sine <= 8'd185;
        10'd436: sine <= 8'd184;
        10'd437: sine <= 8'd183;
        10'd438: sine <= 8'd182;
        10'd439: sine <= 8'd182;
        10'd440: sine <= 8'd181;
        10'd441: sine <= 8'd180;
        10'd442: sine <= 8'd180;
        10'd443: sine <= 8'd179;
        10'd444: sine <= 8'd178;
        10'd445: sine <= 8'd177;
        10'd446: sine <= 8'd177;
        10'd447: sine <= 8'd176;
        10'd448: sine <= 8'd175;
        10'd449: sine <= 8'd175;
        10'd450: sine <= 8'd174;
        10'd451: sine <= 8'd173;
        10'd452: sine <= 8'd172;
        10'd453: sine <= 8'd172;
        10'd454: sine <= 8'd171;
        10'd455: sine <= 8'd170;
        10'd456: sine <= 8'd169;
        10'd457: sine <= 8'd169;
        10'd458: sine <= 8'd168;
        10'd459: sine <= 8'd167;
        10'd460: sine <= 8'd167;
        10'd461: sine <= 8'd166;
        10'd462: sine <= 8'd165;
        10'd463: sine <= 8'd164;
        10'd464: sine <= 8'd164;
        10'd465: sine <= 8'd163;
        10'd466: sine <= 8'd162;
        10'd467: sine <= 8'd161;
        10'd468: sine <= 8'd161;
        10'd469: sine <= 8'd160;
        10'd470: sine <= 8'd159;
        10'd471: sine <= 8'd158;
        10'd472: sine <= 8'd158;
        10'd473: sine <= 8'd157;
        10'd474: sine <= 8'd156;
        10'd475: sine <= 8'd155;
        10'd476: sine <= 8'd154;
        10'd477: sine <= 8'd154;
        10'd478: sine <= 8'd153;
        10'd479: sine <= 8'd152;
        10'd480: sine <= 8'd151;
        10'd481: sine <= 8'd151;
        10'd482: sine <= 8'd150;
        10'd483: sine <= 8'd149;
        10'd484: sine <= 8'd148;
        10'd485: sine <= 8'd148;
        10'd486: sine <= 8'd147;
        10'd487: sine <= 8'd146;
        10'd488: sine <= 8'd145;
        10'd489: sine <= 8'd144;
        10'd490: sine <= 8'd144;
        10'd491: sine <= 8'd143;
        10'd492: sine <= 8'd142;
        10'd493: sine <= 8'd141;
        10'd494: sine <= 8'd141;
        10'd495: sine <= 8'd140;
        10'd496: sine <= 8'd139;
        10'd497: sine <= 8'd138;
        10'd498: sine <= 8'd138;
        10'd499: sine <= 8'd137;
        10'd500: sine <= 8'd136;
        10'd501: sine <= 8'd135;
        10'd502: sine <= 8'd134;
        10'd503: sine <= 8'd134;
        10'd504: sine <= 8'd133;
        10'd505: sine <= 8'd132;
        10'd506: sine <= 8'd131;
        10'd507: sine <= 8'd131;
        10'd508: sine <= 8'd130;
        10'd509: sine <= 8'd129;
        10'd510: sine <= 8'd128;
        10'd511: sine <= 8'd127;
        10'd512: sine <= 8'd127;
        10'd513: sine <= 8'd126;
        10'd514: sine <= 8'd125;
        10'd515: sine <= 8'd124;
        10'd516: sine <= 8'd123;
        10'd517: sine <= 8'd123;
        10'd518: sine <= 8'd122;
        10'd519: sine <= 8'd121;
        10'd520: sine <= 8'd120;
        10'd521: sine <= 8'd120;
        10'd522: sine <= 8'd119;
        10'd523: sine <= 8'd118;
        10'd524: sine <= 8'd117;
        10'd525: sine <= 8'd116;
        10'd526: sine <= 8'd116;
        10'd527: sine <= 8'd115;
        10'd528: sine <= 8'd114;
        10'd529: sine <= 8'd113;
        10'd530: sine <= 8'd113;
        10'd531: sine <= 8'd112;
        10'd532: sine <= 8'd111;
        10'd533: sine <= 8'd110;
        10'd534: sine <= 8'd110;
        10'd535: sine <= 8'd109;
        10'd536: sine <= 8'd108;
        10'd537: sine <= 8'd107;
        10'd538: sine <= 8'd106;
        10'd539: sine <= 8'd106;
        10'd540: sine <= 8'd105;
        10'd541: sine <= 8'd104;
        10'd542: sine <= 8'd103;
        10'd543: sine <= 8'd103;
        10'd544: sine <= 8'd102;
        10'd545: sine <= 8'd101;
        10'd546: sine <= 8'd100;
        10'd547: sine <= 8'd100;
        10'd548: sine <= 8'd99;
        10'd549: sine <= 8'd98;
        10'd550: sine <= 8'd97;
        10'd551: sine <= 8'd96;
        10'd552: sine <= 8'd96;
        10'd553: sine <= 8'd95;
        10'd554: sine <= 8'd94;
        10'd555: sine <= 8'd93;
        10'd556: sine <= 8'd93;
        10'd557: sine <= 8'd92;
        10'd558: sine <= 8'd91;
        10'd559: sine <= 8'd90;
        10'd560: sine <= 8'd90;
        10'd561: sine <= 8'd89;
        10'd562: sine <= 8'd88;
        10'd563: sine <= 8'd87;
        10'd564: sine <= 8'd87;
        10'd565: sine <= 8'd86;
        10'd566: sine <= 8'd85;
        10'd567: sine <= 8'd85;
        10'd568: sine <= 8'd84;
        10'd569: sine <= 8'd83;
        10'd570: sine <= 8'd82;
        10'd571: sine <= 8'd82;
        10'd572: sine <= 8'd81;
        10'd573: sine <= 8'd80;
        10'd574: sine <= 8'd79;
        10'd575: sine <= 8'd79;
        10'd576: sine <= 8'd78;
        10'd577: sine <= 8'd77;
        10'd578: sine <= 8'd77;
        10'd579: sine <= 8'd76;
        10'd580: sine <= 8'd75;
        10'd581: sine <= 8'd74;
        10'd582: sine <= 8'd74;
        10'd583: sine <= 8'd73;
        10'd584: sine <= 8'd72;
        10'd585: sine <= 8'd72;
        10'd586: sine <= 8'd71;
        10'd587: sine <= 8'd70;
        10'd588: sine <= 8'd69;
        10'd589: sine <= 8'd69;
        10'd590: sine <= 8'd68;
        10'd591: sine <= 8'd67;
        10'd592: sine <= 8'd67;
        10'd593: sine <= 8'd66;
        10'd594: sine <= 8'd65;
        10'd595: sine <= 8'd65;
        10'd596: sine <= 8'd64;
        10'd597: sine <= 8'd63;
        10'd598: sine <= 8'd63;
        10'd599: sine <= 8'd62;
        10'd600: sine <= 8'd61;
        10'd601: sine <= 8'd61;
        10'd602: sine <= 8'd60;
        10'd603: sine <= 8'd59;
        10'd604: sine <= 8'd59;
        10'd605: sine <= 8'd58;
        10'd606: sine <= 8'd57;
        10'd607: sine <= 8'd57;
        10'd608: sine <= 8'd56;
        10'd609: sine <= 8'd55;
        10'd610: sine <= 8'd55;
        10'd611: sine <= 8'd54;
        10'd612: sine <= 8'd53;
        10'd613: sine <= 8'd53;
        10'd614: sine <= 8'd52;
        10'd615: sine <= 8'd52;
        10'd616: sine <= 8'd51;
        10'd617: sine <= 8'd50;
        10'd618: sine <= 8'd50;
        10'd619: sine <= 8'd49;
        10'd620: sine <= 8'd48;
        10'd621: sine <= 8'd48;
        10'd622: sine <= 8'd47;
        10'd623: sine <= 8'd47;
        10'd624: sine <= 8'd46;
        10'd625: sine <= 8'd45;
        10'd626: sine <= 8'd45;
        10'd627: sine <= 8'd44;
        10'd628: sine <= 8'd44;
        10'd629: sine <= 8'd43;
        10'd630: sine <= 8'd43;
        10'd631: sine <= 8'd42;
        10'd632: sine <= 8'd41;
        10'd633: sine <= 8'd41;
        10'd634: sine <= 8'd40;
        10'd635: sine <= 8'd40;
        10'd636: sine <= 8'd39;
        10'd637: sine <= 8'd39;
        10'd638: sine <= 8'd38;
        10'd639: sine <= 8'd37;
        10'd640: sine <= 8'd37;
        10'd641: sine <= 8'd36;
        10'd642: sine <= 8'd36;
        10'd643: sine <= 8'd35;
        10'd644: sine <= 8'd35;
        10'd645: sine <= 8'd34;
        10'd646: sine <= 8'd34;
        10'd647: sine <= 8'd33;
        10'd648: sine <= 8'd33;
        10'd649: sine <= 8'd32;
        10'd650: sine <= 8'd32;
        10'd651: sine <= 8'd31;
        10'd652: sine <= 8'd31;
        10'd653: sine <= 8'd30;
        10'd654: sine <= 8'd30;
        10'd655: sine <= 8'd29;
        10'd656: sine <= 8'd29;
        10'd657: sine <= 8'd28;
        10'd658: sine <= 8'd28;
        10'd659: sine <= 8'd27;
        10'd660: sine <= 8'd27;
        10'd661: sine <= 8'd26;
        10'd662: sine <= 8'd26;
        10'd663: sine <= 8'd25;
        10'd664: sine <= 8'd25;
        10'd665: sine <= 8'd24;
        10'd666: sine <= 8'd24;
        10'd667: sine <= 8'd23;
        10'd668: sine <= 8'd23;
        10'd669: sine <= 8'd22;
        10'd670: sine <= 8'd22;
        10'd671: sine <= 8'd22;
        10'd672: sine <= 8'd21;
        10'd673: sine <= 8'd21;
        10'd674: sine <= 8'd20;
        10'd675: sine <= 8'd20;
        10'd676: sine <= 8'd19;
        10'd677: sine <= 8'd19;
        10'd678: sine <= 8'd19;
        10'd679: sine <= 8'd18;
        10'd680: sine <= 8'd18;
        10'd681: sine <= 8'd17;
        10'd682: sine <= 8'd17;
        10'd683: sine <= 8'd17;
        10'd684: sine <= 8'd16;
        10'd685: sine <= 8'd16;
        10'd686: sine <= 8'd15;
        10'd687: sine <= 8'd15;
        10'd688: sine <= 8'd15;
        10'd689: sine <= 8'd14;
        10'd690: sine <= 8'd14;
        10'd691: sine <= 8'd14;
        10'd692: sine <= 8'd13;
        10'd693: sine <= 8'd13;
        10'd694: sine <= 8'd13;
        10'd695: sine <= 8'd12;
        10'd696: sine <= 8'd12;
        10'd697: sine <= 8'd12;
        10'd698: sine <= 8'd11;
        10'd699: sine <= 8'd11;
        10'd700: sine <= 8'd11;
        10'd701: sine <= 8'd10;
        10'd702: sine <= 8'd10;
        10'd703: sine <= 8'd10;
        10'd704: sine <= 8'd9;
        10'd705: sine <= 8'd9;
        10'd706: sine <= 8'd9;
        10'd707: sine <= 8'd9;
        10'd708: sine <= 8'd8;
        10'd709: sine <= 8'd8;
        10'd710: sine <= 8'd8;
        10'd711: sine <= 8'd8;
        10'd712: sine <= 8'd7;
        10'd713: sine <= 8'd7;
        10'd714: sine <= 8'd7;
        10'd715: sine <= 8'd6;
        10'd716: sine <= 8'd6;
        10'd717: sine <= 8'd6;
        10'd718: sine <= 8'd6;
        10'd719: sine <= 8'd6;
        10'd720: sine <= 8'd5;
        10'd721: sine <= 8'd5;
        10'd722: sine <= 8'd5;
        10'd723: sine <= 8'd5;
        10'd724: sine <= 8'd4;
        10'd725: sine <= 8'd4;
        10'd726: sine <= 8'd4;
        10'd727: sine <= 8'd4;
        10'd728: sine <= 8'd4;
        10'd729: sine <= 8'd3;
        10'd730: sine <= 8'd3;
        10'd731: sine <= 8'd3;
        10'd732: sine <= 8'd3;
        10'd733: sine <= 8'd3;
        10'd734: sine <= 8'd3;
        10'd735: sine <= 8'd2;
        10'd736: sine <= 8'd2;
        10'd737: sine <= 8'd2;
        10'd738: sine <= 8'd2;
        10'd739: sine <= 8'd2;
        10'd740: sine <= 8'd2;
        10'd741: sine <= 8'd2;
        10'd742: sine <= 8'd2;
        10'd743: sine <= 8'd1;
        10'd744: sine <= 8'd1;
        10'd745: sine <= 8'd1;
        10'd746: sine <= 8'd1;
        10'd747: sine <= 8'd1;
        10'd748: sine <= 8'd1;
        10'd749: sine <= 8'd1;
        10'd750: sine <= 8'd1;
        10'd751: sine <= 8'd1;
        10'd752: sine <= 8'd1;
        10'd753: sine <= 8'd0;
        10'd754: sine <= 8'd0;
        10'd755: sine <= 8'd0;
        10'd756: sine <= 8'd0;
        10'd757: sine <= 8'd0;
        10'd758: sine <= 8'd0;
        10'd759: sine <= 8'd0;
        10'd760: sine <= 8'd0;
        10'd761: sine <= 8'd0;
        10'd762: sine <= 8'd0;
        10'd763: sine <= 8'd0;
        10'd764: sine <= 8'd0;
        10'd765: sine <= 8'd0;
        10'd766: sine <= 8'd0;
        10'd767: sine <= 8'd0;
        10'd768: sine <= 8'd0;
        10'd769: sine <= 8'd0;
        10'd770: sine <= 8'd0;
        10'd771: sine <= 8'd0;
        10'd772: sine <= 8'd0;
        10'd773: sine <= 8'd0;
        10'd774: sine <= 8'd0;
        10'd775: sine <= 8'd0;
        10'd776: sine <= 8'd0;
        10'd777: sine <= 8'd0;
        10'd778: sine <= 8'd0;
        10'd779: sine <= 8'd0;
        10'd780: sine <= 8'd0;
        10'd781: sine <= 8'd0;
        10'd782: sine <= 8'd1;
        10'd783: sine <= 8'd1;
        10'd784: sine <= 8'd1;
        10'd785: sine <= 8'd1;
        10'd786: sine <= 8'd1;
        10'd787: sine <= 8'd1;
        10'd788: sine <= 8'd1;
        10'd789: sine <= 8'd1;
        10'd790: sine <= 8'd1;
        10'd791: sine <= 8'd1;
        10'd792: sine <= 8'd1;
        10'd793: sine <= 8'd2;
        10'd794: sine <= 8'd2;
        10'd795: sine <= 8'd2;
        10'd796: sine <= 8'd2;
        10'd797: sine <= 8'd2;
        10'd798: sine <= 8'd2;
        10'd799: sine <= 8'd2;
        10'd800: sine <= 8'd3;
        10'd801: sine <= 8'd3;
        10'd802: sine <= 8'd3;
        10'd803: sine <= 8'd3;
        10'd804: sine <= 8'd3;
        10'd805: sine <= 8'd3;
        10'd806: sine <= 8'd4;
        10'd807: sine <= 8'd4;
        10'd808: sine <= 8'd4;
        10'd809: sine <= 8'd4;
        10'd810: sine <= 8'd4;
        10'd811: sine <= 8'd5;
        10'd812: sine <= 8'd5;
        10'd813: sine <= 8'd5;
        10'd814: sine <= 8'd5;
        10'd815: sine <= 8'd5;
        10'd816: sine <= 8'd6;
        10'd817: sine <= 8'd6;
        10'd818: sine <= 8'd6;
        10'd819: sine <= 8'd6;
        10'd820: sine <= 8'd7;
        10'd821: sine <= 8'd7;
        10'd822: sine <= 8'd7;
        10'd823: sine <= 8'd7;
        10'd824: sine <= 8'd8;
        10'd825: sine <= 8'd8;
        10'd826: sine <= 8'd8;
        10'd827: sine <= 8'd8;
        10'd828: sine <= 8'd9;
        10'd829: sine <= 8'd9;
        10'd830: sine <= 8'd9;
        10'd831: sine <= 8'd10;
        10'd832: sine <= 8'd10;
        10'd833: sine <= 8'd10;
        10'd834: sine <= 8'd11;
        10'd835: sine <= 8'd11;
        10'd836: sine <= 8'd11;
        10'd837: sine <= 8'd11;
        10'd838: sine <= 8'd12;
        10'd839: sine <= 8'd12;
        10'd840: sine <= 8'd12;
        10'd841: sine <= 8'd13;
        10'd842: sine <= 8'd13;
        10'd843: sine <= 8'd13;
        10'd844: sine <= 8'd14;
        10'd845: sine <= 8'd14;
        10'd846: sine <= 8'd15;
        10'd847: sine <= 8'd15;
        10'd848: sine <= 8'd15;
        10'd849: sine <= 8'd16;
        10'd850: sine <= 8'd16;
        10'd851: sine <= 8'd16;
        10'd852: sine <= 8'd17;
        10'd853: sine <= 8'd17;
        10'd854: sine <= 8'd18;
        10'd855: sine <= 8'd18;
        10'd856: sine <= 8'd18;
        10'd857: sine <= 8'd19;
        10'd858: sine <= 8'd19;
        10'd859: sine <= 8'd20;
        10'd860: sine <= 8'd20;
        10'd861: sine <= 8'd20;
        10'd862: sine <= 8'd21;
        10'd863: sine <= 8'd21;
        10'd864: sine <= 8'd22;
        10'd865: sine <= 8'd22;
        10'd866: sine <= 8'd23;
        10'd867: sine <= 8'd23;
        10'd868: sine <= 8'd24;
        10'd869: sine <= 8'd24;
        10'd870: sine <= 8'd24;
        10'd871: sine <= 8'd25;
        10'd872: sine <= 8'd25;
        10'd873: sine <= 8'd26;
        10'd874: sine <= 8'd26;
        10'd875: sine <= 8'd27;
        10'd876: sine <= 8'd27;
        10'd877: sine <= 8'd28;
        10'd878: sine <= 8'd28;
        10'd879: sine <= 8'd29;
        10'd880: sine <= 8'd29;
        10'd881: sine <= 8'd30;
        10'd882: sine <= 8'd30;
        10'd883: sine <= 8'd31;
        10'd884: sine <= 8'd31;
        10'd885: sine <= 8'd32;
        10'd886: sine <= 8'd32;
        10'd887: sine <= 8'd33;
        10'd888: sine <= 8'd33;
        10'd889: sine <= 8'd34;
        10'd890: sine <= 8'd34;
        10'd891: sine <= 8'd35;
        10'd892: sine <= 8'd35;
        10'd893: sine <= 8'd36;
        10'd894: sine <= 8'd37;
        10'd895: sine <= 8'd37;
        10'd896: sine <= 8'd38;
        10'd897: sine <= 8'd38;
        10'd898: sine <= 8'd39;
        10'd899: sine <= 8'd39;
        10'd900: sine <= 8'd40;
        10'd901: sine <= 8'd40;
        10'd902: sine <= 8'd41;
        10'd903: sine <= 8'd42;
        10'd904: sine <= 8'd42;
        10'd905: sine <= 8'd43;
        10'd906: sine <= 8'd43;
        10'd907: sine <= 8'd44;
        10'd908: sine <= 8'd45;
        10'd909: sine <= 8'd45;
        10'd910: sine <= 8'd46;
        10'd911: sine <= 8'd46;
        10'd912: sine <= 8'd47;
        10'd913: sine <= 8'd48;
        10'd914: sine <= 8'd48;
        10'd915: sine <= 8'd49;
        10'd916: sine <= 8'd49;
        10'd917: sine <= 8'd50;
        10'd918: sine <= 8'd51;
        10'd919: sine <= 8'd51;
        10'd920: sine <= 8'd52;
        10'd921: sine <= 8'd53;
        10'd922: sine <= 8'd53;
        10'd923: sine <= 8'd54;
        10'd924: sine <= 8'd54;
        10'd925: sine <= 8'd55;
        10'd926: sine <= 8'd56;
        10'd927: sine <= 8'd56;
        10'd928: sine <= 8'd57;
        10'd929: sine <= 8'd58;
        10'd930: sine <= 8'd58;
        10'd931: sine <= 8'd59;
        10'd932: sine <= 8'd60;
        10'd933: sine <= 8'd60;
        10'd934: sine <= 8'd61;
        10'd935: sine <= 8'd62;
        10'd936: sine <= 8'd62;
        10'd937: sine <= 8'd63;
        10'd938: sine <= 8'd64;
        10'd939: sine <= 8'd64;
        10'd940: sine <= 8'd65;
        10'd941: sine <= 8'd66;
        10'd942: sine <= 8'd66;
        10'd943: sine <= 8'd67;
        10'd944: sine <= 8'd68;
        10'd945: sine <= 8'd68;
        10'd946: sine <= 8'd69;
        10'd947: sine <= 8'd70;
        10'd948: sine <= 8'd71;
        10'd949: sine <= 8'd71;
        10'd950: sine <= 8'd72;
        10'd951: sine <= 8'd73;
        10'd952: sine <= 8'd73;
        10'd953: sine <= 8'd74;
        10'd954: sine <= 8'd75;
        10'd955: sine <= 8'd75;
        10'd956: sine <= 8'd76;
        10'd957: sine <= 8'd77;
        10'd958: sine <= 8'd78;
        10'd959: sine <= 8'd78;
        10'd960: sine <= 8'd79;
        10'd961: sine <= 8'd80;
        10'd962: sine <= 8'd81;
        10'd963: sine <= 8'd81;
        10'd964: sine <= 8'd82;
        10'd965: sine <= 8'd83;
        10'd966: sine <= 8'd83;
        10'd967: sine <= 8'd84;
        10'd968: sine <= 8'd85;
        10'd969: sine <= 8'd86;
        10'd970: sine <= 8'd86;
        10'd971: sine <= 8'd87;
        10'd972: sine <= 8'd88;
        10'd973: sine <= 8'd89;
        10'd974: sine <= 8'd89;
        10'd975: sine <= 8'd90;
        10'd976: sine <= 8'd91;
        10'd977: sine <= 8'd92;
        10'd978: sine <= 8'd92;
        10'd979: sine <= 8'd93;
        10'd980: sine <= 8'd94;
        10'd981: sine <= 8'd95;
        10'd982: sine <= 8'd95;
        10'd983: sine <= 8'd96;
        10'd984: sine <= 8'd97;
        10'd985: sine <= 8'd98;
        10'd986: sine <= 8'd98;
        10'd987: sine <= 8'd99;
        10'd988: sine <= 8'd100;
        10'd989: sine <= 8'd101;
        10'd990: sine <= 8'd101;
        10'd991: sine <= 8'd102;
        10'd992: sine <= 8'd103;
        10'd993: sine <= 8'd104;
        10'd994: sine <= 8'd104;
        10'd995: sine <= 8'd105;
        10'd996: sine <= 8'd106;
        10'd997: sine <= 8'd107;
        10'd998: sine <= 8'd108;
        10'd999: sine <= 8'd108;
        10'd1000: sine <= 8'd109;
        10'd1001: sine <= 8'd110;
        10'd1002: sine <= 8'd111;
        10'd1003: sine <= 8'd111;
        10'd1004: sine <= 8'd112;
        10'd1005: sine <= 8'd113;
        10'd1006: sine <= 8'd114;
        10'd1007: sine <= 8'd115;
        10'd1008: sine <= 8'd115;
        10'd1009: sine <= 8'd116;
        10'd1010: sine <= 8'd117;
        10'd1011: sine <= 8'd118;
        10'd1012: sine <= 8'd118;
        10'd1013: sine <= 8'd119;
        10'd1014: sine <= 8'd120;
        10'd1015: sine <= 8'd121;
        10'd1016: sine <= 8'd122;
        10'd1017: sine <= 8'd122;
        10'd1018: sine <= 8'd123;
        10'd1019: sine <= 8'd124;
        10'd1020: sine <= 8'd125;
        10'd1021: sine <= 8'd125;
        10'd1022: sine <= 8'd126;
        10'd1023: sine <= 8'd127;
    endcase
end
endmodule
